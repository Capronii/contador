library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 13;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is
  
  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI	 : std_logic_vector(3 downto 0) := "0100";
  constant STA	 : std_logic_vector(3 downto 0) := "0101";
  constant JMP : std_logic_vector(3 downto 0) := "0110";
  constant JEQ : std_logic_vector(3 downto 0) := "0111";
  constant CEQ : std_logic_vector(3 downto 0) := "1000";
  constant JSR : std_logic_vector(3 downto 0) := "1001";
  constant RET : std_logic_vector(3 downto 0) := "1010";
  constant GT : std_logic_vector(3 downto 0) := "1011";
  constant JGT : std_logic_vector(3 downto 0) := "1100";


  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
      -- Palavra de Controle = SelMUX, Habilita_A, Reset_A, Operacao_ULA
      -- Inicializa os endereços:
tmp(0) := NOP & '0' & x"00";	-- NOP 
tmp(1) := LDI & '0' & x"00";	-- LDI $0    	#Início do Setup
tmp(2) := STA & '1' & x"20";	-- STA @288    	#Zerando hexas
tmp(3) := STA & '1' & x"21";	-- STA @289
tmp(4) := STA & '1' & x"22";	-- STA @290
tmp(5) := STA & '1' & x"23";	-- STA @291
tmp(6) := STA & '1' & x"24";	-- STA @292
tmp(7) := STA & '1' & x"25";	-- STA @293
tmp(8) := STA & '1' & x"00";	-- STA @256    	#Zerando leds
tmp(9) := STA & '1' & x"01";	-- STA @257
tmp(10) := STA & '1' & x"02";	-- STA @258
tmp(11) := STA & '0' & x"00";	-- STA @0    	#Armazenando 0 em unidade, dezena, centena, etc
tmp(12) := STA & '0' & x"01";	-- STA @1
tmp(13) := STA & '0' & x"02";	-- STA @2
tmp(14) := STA & '0' & x"03";	-- STA @3
tmp(15) := STA & '0' & x"04";	-- STA @4
tmp(16) := STA & '0' & x"05";	-- STA @5
tmp(17) := STA & '0' & x"06";	-- STA @6    	#Constante de comparacao (0)
tmp(18) := STA & '0' & x"0F";	-- STA @15   	#Flag que para contagem
tmp(19) := STA & '1' & x"FE";	-- STA @510
tmp(20) := STA & '1' & x"FF";	-- STA @511
tmp(21) := STA & '1' & x"FD";	-- STA @509
tmp(22) := LDI & '0' & x"01";	-- LDI $1
tmp(23) := STA & '0' & x"07";	-- STA @7    	#Constante de Incremento (1)
tmp(24) := LDI & '0' & x"0A";	-- LDI $10
tmp(25) := STA & '0' & x"08";	-- STA @8    	#Constante de limite no display (10)
tmp(26) := LDI & '0' & x"00";	-- LDI $0
tmp(27) := STA & '0' & x"09";	-- STA @9    	#Limite de contagem em unidade, dezena, centena, etc
tmp(28) := STA & '0' & x"0A";	-- STA @10  
tmp(29) := STA & '0' & x"0B";	-- STA @11
tmp(30) := STA & '0' & x"0C";	-- STA @12
tmp(31) := STA & '0' & x"0D";	-- STA @13
tmp(32) := STA & '0' & x"0E";	-- STA @14
tmp(33) := LDI & '0' & x"0B";	-- LDI $11
tmp(34) := STA & '0' & x"10";	-- STA @16   	#Constante de limite de contagem (11)
tmp(35) := LDI & '0' & x"0C";	-- LDI $12
tmp(36) := STA & '0' & x"11";	-- STA @17   	#Constante de limite de contagem (12)
tmp(37) := LDI & '0' & x"0D";	-- LDI $13
tmp(38) := STA & '0' & x"12";	-- STA @18   	#Constante de limite de contagem (13)
tmp(39) := LDI & '0' & x"0E";	-- LDI $14
tmp(40) := STA & '0' & x"13";	-- STA @19   	#Constante de limite de contagem (14)
tmp(41) := LDI & '0' & x"0F";	-- LDI $15 
tmp(42) := STA & '0' & x"14";	-- STA @20   	#Constante de limite de contagem (15)
tmp(43) := LDI & '0' & x"00";	-- LDI $0
tmp(44) := STA & '0' & x"15";	-- STA @21   	#Constante de limite de contagem (0)
tmp(45) := NOP & '0' & x"00";	-- NOP  	#Loop principal
tmp(46) := LDA & '1' & x"61";	-- LDA @353 	# Le o valor de KEY1
tmp(47) := CEQ & '0' & x"06";	-- CEQ @6 	# Compara o valor de KEY1 com 0
tmp(48) := JEQ & '0' & x"2D";	-- JEQ @INICIOLOOP 	# Se for igual a 0, fica no aguardo para quando for 1
tmp(49) := JSR & '0' & x"48";	-- JSR @CONFIGLIMITE 	# Se for diferente de 0, entra na sub rotina de configuracao de Limite
tmp(50) := LDA & '0' & x"06";	-- LDA @6 	#Carrega 0 no acumulador
tmp(51) := STA & '1' & x"20";	-- STA @288 	# Zera o HEX1
tmp(52) := STA & '1' & x"21";	-- STA @289 	# Zera o HEX2
tmp(53) := STA & '1' & x"22";	-- STA @290 	# Zera o HEX3
tmp(54) := STA & '1' & x"23";	-- STA @291 	# Zera o HEX4
tmp(55) := STA & '1' & x"24";	-- STA @292 	# Zera o HEX5
tmp(56) := STA & '1' & x"25";	-- STA @293 	# Zera o HEX6
tmp(57) := STA & '1' & x"00";	-- STA @256 	# Zera os LEDS(7~0)
tmp(58) := STA & '1' & x"02";	-- STA @258 	# Zera os LED(9)
tmp(59) := STA & '1' & x"01";	-- STA @257 	# Zera os LED(8) 
tmp(60) := NOP & '0' & x"00";	-- NOP  	# Incrementa ate chegar no limite de contagem
tmp(61) := LDA & '1' & x"60";	-- LDA @352 	# Le o valor de KEY0
tmp(62) := CEQ & '0' & x"06";	-- CEQ @6   	# Compara o valor de KEY0 com 0
tmp(63) := JEQ & '0' & x"41";	-- JEQ @PULA1 	# Se for igual a 0, nao incrementa e atualiza os displays
tmp(64) := JSR & '1' & x"2B";	-- JSR @INCREMENTA 	# Se for diferente de 0, entra na sub rotina de incremento
tmp(65) := NOP & '0' & x"00";	-- NOP 
tmp(66) := JSR & '1' & x"68";	-- JSR @ATUALIZA 	# Atualiza os displays
tmp(67) := JSR & '1' & x"76";	-- JSR @CHECALIMITE 	# Checa pra ver se passou do limite setado
tmp(68) := LDA & '0' & x"0F";	-- LDA @15 	# Le o valor da flag de inibir contagem
tmp(69) := CEQ & '0' & x"06";	-- CEQ @6 	# Compara com 0 a flag (flag com valor 1 -> ativa, flag com valor 0 -> desativada)
tmp(70) := JEQ & '0' & x"3C";	-- JEQ @INCREMENTADOR 	#Se a flag for 0, pode continuar incrementando
tmp(71) := JMP & '1' & x"99";	-- JMP @TRAVA 	# Se for 1, trava a contagem
tmp(72) := NOP & '0' & x"00";	-- NOP  	#Rotina de configuracao de limite
tmp(73) := LDI & '0' & x"01";	-- LDI $1 	# Carrega o valor 1
tmp(74) := STA & '1' & x"00";	-- STA @256 	# Bota no endereco dos LEDS(7-0)
tmp(75) := STA & '1' & x"FE";	-- STA @510 	#Limpa a leitura de KEY1
tmp(76) := NOP & '0' & x"00";	-- NOP 
tmp(77) := LDA & '1' & x"40";	-- LDA @320 	#Le o valor das chaves SW(7~0)
tmp(78) := CEQ & '0' & x"08";	-- CEQ @8 	#Compara com 10
tmp(79) := JEQ & '1' & x"A0";	-- JEQ @DISPLAYATUALIZADO0 	#Se for 10, atualiza o display e vai para a proxima configuracao
tmp(80) := CEQ & '0' & x"10";	-- CEQ @16 	#Compara com 11 
tmp(81) := JEQ & '1' & x"A0";	-- JEQ @DISPLAYATUALIZADO0 	#Se for 11, atualiza o display e vai para a proxima configuracao
tmp(82) := CEQ & '0' & x"11";	-- CEQ @17 	#Compara com 12 
tmp(83) := JEQ & '1' & x"A0";	-- JEQ @DISPLAYATUALIZADO0 	#Se for 12, atualiza o display e vai para a proxima configuracao
tmp(84) := CEQ & '0' & x"12";	-- CEQ @18 	#Compara com 13
tmp(85) := JEQ & '1' & x"A0";	-- JEQ @DISPLAYATUALIZADO0 	#Se for 13, atualiza o display e vai para a proxima configuracao
tmp(86) := CEQ & '0' & x"13";	-- CEQ @19 	#Compara com 14
tmp(87) := JEQ & '1' & x"A0";	-- JEQ @DISPLAYATUALIZADO0 	#Se for 14, atualiza o display e vai para a proxima configuracao
tmp(88) := CEQ & '0' & x"14";	-- CEQ @20 	#Compara com 15
tmp(89) := JEQ & '1' & x"A0";	-- JEQ @DISPLAYATUALIZADO0 	#Se for 15, atualiza o display e vai para a proxima configuracao
tmp(90) := NOP & '0' & x"00";	-- NOP 
tmp(91) := STA & '1' & x"20";	-- STA @288 	# Hex 0
tmp(92) := LDA & '1' & x"61";	-- LDA @353 	# Le KEY1
tmp(93) := CEQ & '0' & x"06";	-- CEQ @6 	#Compara KEY1 com 0
tmp(94) := JEQ & '0' & x"4C";	-- JEQ @ESPERAUNIDADE  	#Se for 0, ou seja, nao esta apertado, espera ate apertar
tmp(95) := STA & '1' & x"FE";	-- STA @510 	#Limpa a leitura de KEY1
tmp(96) := LDA & '1' & x"40";	-- LDA @320 	#Le o valor das chaves SW(7~0)
tmp(97) := CEQ & '0' & x"08";	-- CEQ @8 	#Compara com 10
tmp(98) := JEQ & '1' & x"B2";	-- JEQ @VALORATUALIZADO0 	#Se for 10, atualiza o valor e vai para a proxima configuracao
tmp(99) := CEQ & '0' & x"10";	-- CEQ @16 	#Compara com 11
tmp(100) := JEQ & '1' & x"B2";	-- JEQ @VALORATUALIZADO0 	#Se for 11, atualiza o valor e vai para a proxima configuracao
tmp(101) := CEQ & '0' & x"11";	-- CEQ @17 	#Compara com 12
tmp(102) := JEQ & '1' & x"B2";	-- JEQ @VALORATUALIZADO0 	#Se for 12, atualiza o valor e vai para a proxima configuracao
tmp(103) := CEQ & '0' & x"12";	-- CEQ @18 	#Compara com 13
tmp(104) := JEQ & '1' & x"B2";	-- JEQ @VALORATUALIZADO0 	#Se for 13, atualiza o valor e vai para a proxima configuracao
tmp(105) := CEQ & '0' & x"13";	-- CEQ @19 	#Compara com 14
tmp(106) := JEQ & '1' & x"B2";	-- JEQ @VALORATUALIZADO0 	#Se for 14, atualiza o valor e vai para a proxima configuracao
tmp(107) := CEQ & '0' & x"14";	-- CEQ @20 	#Compara com 15
tmp(108) := JEQ & '1' & x"B2";	-- JEQ @VALORATUALIZADO0 	#Se for 15, atualiza o valor e vai para a proxima configuracao
tmp(109) := NOP & '0' & x"00";	-- NOP 
tmp(110) := STA & '0' & x"09";	-- STA @9   	#Armazena o valor das chaves no limite das unidades
tmp(111) := NOP & '0' & x"00";	-- NOP 
tmp(112) := LDI & '0' & x"04";	-- LDI $4 	#Carrega o valor 4
tmp(113) := STA & '1' & x"00";	-- STA @256 	# Bota o valor nos LEDS
tmp(114) := LDA & '1' & x"40";	-- LDA @320 	#Le o valor das chaves SW(7~0)
tmp(115) := CEQ & '0' & x"08";	-- CEQ @8 	#Compara com 10
tmp(116) := JEQ & '1' & x"A3";	-- JEQ @DISPLAYATUALIZADO1 	#Se for 10, atualiza o display e vai para a proxima configuracao
tmp(117) := CEQ & '0' & x"10";	-- CEQ @16 	#Compara com 11
tmp(118) := JEQ & '1' & x"A3";	-- JEQ @DISPLAYATUALIZADO1 	#Se for 11, atualiza o display e vai para a proxima configuracao
tmp(119) := CEQ & '0' & x"11";	-- CEQ @17 	#Compara com 12
tmp(120) := JEQ & '1' & x"A3";	-- JEQ @DISPLAYATUALIZADO1 	#Se for 12, atualiza o display e vai para a proxima configuracao
tmp(121) := CEQ & '0' & x"12";	-- CEQ @18 	#Compara com 13
tmp(122) := JEQ & '1' & x"A3";	-- JEQ @DISPLAYATUALIZADO1 	#Se for 13, atualiza o display e vai para a proxima configuracao
tmp(123) := CEQ & '0' & x"13";	-- CEQ @19 	#Compara com 14
tmp(124) := JEQ & '1' & x"A3";	-- JEQ @DISPLAYATUALIZADO1 	#Se for 14, atualiza o display e vai para a proxima configuracao
tmp(125) := CEQ & '0' & x"14";	-- CEQ @20 	#Compara com 15
tmp(126) := JEQ & '1' & x"A3";	-- JEQ @DISPLAYATUALIZADO1 	#Se for 15, atualiza o display e vai para a proxima configuracao
tmp(127) := NOP & '0' & x"00";	-- NOP 
tmp(128) := STA & '1' & x"21";	-- STA @289 	# Hex 1
tmp(129) := LDA & '1' & x"61";	-- LDA @353 	#Le o valor de KEY1 novamente
tmp(130) := CEQ & '0' & x"06";	-- CEQ @6 	#Compara com 0 o valor de KEY1 
tmp(131) := JEQ & '0' & x"6F";	-- JEQ @ESPERADEZENA 	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(132) := STA & '1' & x"FE";	-- STA @510 	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(133) := LDA & '1' & x"40";	-- LDA @320 	#Le o valor das chaves SW(7~0)
tmp(134) := CEQ & '0' & x"08";	-- CEQ @8 	#Compara com 10
tmp(135) := JEQ & '1' & x"B5";	-- JEQ @VALORATUALIZADO1  	#Se for 10, atualiza o valor e vai para a proxima configuracao
tmp(136) := CEQ & '0' & x"10";	-- CEQ @16 	#Compara com 11
tmp(137) := JEQ & '1' & x"B5";	-- JEQ @VALORATUALIZADO1 	#Se for 11, atualiza o valor e vai para a proxima configuracao
tmp(138) := CEQ & '0' & x"11";	-- CEQ @17 	#Compara com 12
tmp(139) := JEQ & '1' & x"B5";	-- JEQ @VALORATUALIZADO1 	#Se for 12, atualiza o valor e vai para a proxima configuracao
tmp(140) := CEQ & '0' & x"12";	-- CEQ @18 	#Compara com 13
tmp(141) := JEQ & '1' & x"B5";	-- JEQ @VALORATUALIZADO1 	#Se for 13, atualiza o valor e vai para a proxima configuracao
tmp(142) := CEQ & '0' & x"13";	-- CEQ @19 	#Compara com 14
tmp(143) := JEQ & '1' & x"B5";	-- JEQ @VALORATUALIZADO1 	#Se for 14, atualiza o valor e vai para a proxima configuracao
tmp(144) := CEQ & '0' & x"14";	-- CEQ @20 	#Compara com 15
tmp(145) := JEQ & '1' & x"B5";	-- JEQ @VALORATUALIZADO1 	#Se for 15, atualiza o valor e vai para a proxima configuracao
tmp(146) := NOP & '0' & x"00";	-- NOP 
tmp(147) := STA & '0' & x"0A";	-- STA @10 	#Armazena o valor das chaves no limte das dezenas
tmp(148) := NOP & '0' & x"00";	-- NOP 
tmp(149) := LDI & '0' & x"10";	-- LDI $16 	# Carrega o valor 16 no acumulador
tmp(150) := STA & '1' & x"00";	-- STA @256 	# Bota o valor nos LEDS
tmp(151) := LDA & '1' & x"40";	-- LDA @320 	#Le o valor das chaves SW(7~0)
tmp(152) := CEQ & '0' & x"08";	-- CEQ @8 	#Compara com 10
tmp(153) := JEQ & '1' & x"A6";	-- JEQ @DISPLAYATUALIZADO2 	#Se for 10, atualiza o display e vai para a proxima configuracao
tmp(154) := CEQ & '0' & x"10";	-- CEQ @16 	#Compara com 11
tmp(155) := JEQ & '1' & x"A6";	-- JEQ @DISPLAYATUALIZADO2 	#Se for 11, atualiza o display e vai para a proxima configuracao
tmp(156) := CEQ & '0' & x"11";	-- CEQ @17 	#Compara com 12
tmp(157) := JEQ & '1' & x"A6";	-- JEQ @DISPLAYATUALIZADO2 	#Se for 12, atualiza o display e vai para a proxima configuracao
tmp(158) := CEQ & '0' & x"12";	-- CEQ @18 	#Compara com 13
tmp(159) := JEQ & '1' & x"A6";	-- JEQ @DISPLAYATUALIZADO2 	#Se for 13, atualiza o display e vai para a proxima configuracao
tmp(160) := CEQ & '0' & x"13";	-- CEQ @19 	#Compara com 14
tmp(161) := JEQ & '1' & x"A6";	-- JEQ @DISPLAYATUALIZADO2 	#Se for 14, atualiza o display e vai para a proxima configuracao
tmp(162) := CEQ & '0' & x"14";	-- CEQ @20 	#Compara com 15
tmp(163) := JEQ & '1' & x"A6";	-- JEQ @DISPLAYATUALIZADO2 	#Se for 15, atualiza o display e vai para a proxima configuracao
tmp(164) := NOP & '0' & x"00";	-- NOP 
tmp(165) := STA & '1' & x"22";	-- STA @290 	# Hex 2
tmp(166) := LDA & '1' & x"61";	-- LDA @353 	#Le o valor de KEY1 novamente
tmp(167) := CEQ & '0' & x"06";	-- CEQ @6 	#Compara com 0 o valor de KEY1 
tmp(168) := JEQ & '0' & x"94";	-- JEQ @ESPERACENTENA 	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(169) := STA & '1' & x"FE";	-- STA @510 	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(170) := LDA & '1' & x"40";	-- LDA @320 	#Le o valor das chaves SW(7~0)
tmp(171) := CEQ & '0' & x"08";	-- CEQ @8 	#Compara com 10
tmp(172) := JEQ & '1' & x"B8";	-- JEQ @VALORATUALIZADO2 	#Se for 10, atualiza o valor e vai para a proxima configuracao
tmp(173) := CEQ & '0' & x"10";	-- CEQ @16 	#Compara com 11
tmp(174) := JEQ & '1' & x"B8";	-- JEQ @VALORATUALIZADO2 	#Se for 11, atualiza o valor e vai para a proxima configuracao
tmp(175) := CEQ & '0' & x"11";	-- CEQ @17 	#Compara com 12
tmp(176) := JEQ & '1' & x"B8";	-- JEQ @VALORATUALIZADO2 	#Se for 12, atualiza o valor e vai para a proxima configuracao
tmp(177) := CEQ & '0' & x"12";	-- CEQ @18 	#Compara com 13
tmp(178) := JEQ & '1' & x"B8";	-- JEQ @VALORATUALIZADO2 	#Se for 13, atualiza o valor e vai para a proxima configuracao
tmp(179) := CEQ & '0' & x"13";	-- CEQ @19 	#Compara com 14
tmp(180) := JEQ & '1' & x"B8";	-- JEQ @VALORATUALIZADO2   	#Se for 14, atualiza o valor e vai para a proxima configuracao
tmp(181) := CEQ & '0' & x"14";	-- CEQ @20 	#Compara com 15
tmp(182) := JEQ & '1' & x"B8";	-- JEQ @VALORATUALIZADO2 	#Se for 15, atualiza o valor e vai para a proxima configuracao
tmp(183) := NOP & '0' & x"00";	-- NOP 
tmp(184) := STA & '0' & x"0B";	-- STA @11 	#Armazena o valor das chaves no limite das centenas
tmp(185) := NOP & '0' & x"00";	-- NOP 
tmp(186) := LDI & '0' & x"20";	-- LDI $32 	# Carrega o valor 32 no acumulador
tmp(187) := STA & '1' & x"00";	-- STA @256 	# Bota o valor nos LEDS
tmp(188) := LDA & '1' & x"40";	-- LDA @320 	#Le o valor das chaves SW(7~0)
tmp(189) := CEQ & '0' & x"08";	-- CEQ @8 	#Compara com 10
tmp(190) := JEQ & '1' & x"A9";	-- JEQ @DISPLAYATUALIZADO3 	#Se for 10, atualiza o display e vai para a proxima configuracao
tmp(191) := CEQ & '0' & x"10";	-- CEQ @16 	#Compara com 11
tmp(192) := JEQ & '1' & x"A9";	-- JEQ @DISPLAYATUALIZADO3 	#Se for 11, atualiza o display e vai para a proxima configuracao
tmp(193) := CEQ & '0' & x"11";	-- CEQ @17 	#Compara com 12
tmp(194) := JEQ & '1' & x"A9";	-- JEQ @DISPLAYATUALIZADO3 	#Se for 12, atualiza o display e vai para a proxima configuracao
tmp(195) := CEQ & '0' & x"12";	-- CEQ @18 	#Compara com 13
tmp(196) := JEQ & '1' & x"A9";	-- JEQ @DISPLAYATUALIZADO3 	#Se for 13, atualiza o display e vai para a proxima configuracao
tmp(197) := CEQ & '0' & x"13";	-- CEQ @19 	#Compara com 14
tmp(198) := JEQ & '1' & x"A9";	-- JEQ @DISPLAYATUALIZADO3 	#Se for 14, atualiza o display e vai para a proxima configuracao
tmp(199) := CEQ & '0' & x"14";	-- CEQ @20 	#Compara com 15
tmp(200) := JEQ & '1' & x"A9";	-- JEQ @DISPLAYATUALIZADO3 	#Se for 15, atualiza o display e vai para a proxima configuracao
tmp(201) := NOP & '0' & x"00";	-- NOP 
tmp(202) := STA & '1' & x"23";	-- STA @291 	# Hex 3
tmp(203) := LDA & '1' & x"61";	-- LDA @353 	#Le o valor de KEY1 novamente
tmp(204) := CEQ & '0' & x"06";	-- CEQ @6 	#Compara com 0 o valor de KEY1
tmp(205) := JEQ & '0' & x"B9";	-- JEQ @ESPERAUNIDADEMILHAR 	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(206) := STA & '1' & x"FE";	-- STA @510 	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(207) := LDA & '1' & x"40";	-- LDA @320 	#Le o valor das chaves SW(7~0)
tmp(208) := CEQ & '0' & x"08";	-- CEQ @8 	#Compara com 10
tmp(209) := JEQ & '1' & x"BB";	-- JEQ @VALORATUALIZADO3 	#Se for 10, atualiza o valor e vai para a proxima configuracao
tmp(210) := CEQ & '0' & x"10";	-- CEQ @16 	#Compara com 11
tmp(211) := JEQ & '1' & x"BB";	-- JEQ @VALORATUALIZADO3 	#Se for 11, atualiza o valor e vai para a proxima configuracao
tmp(212) := CEQ & '0' & x"11";	-- CEQ @17 	#Compara com 12
tmp(213) := JEQ & '1' & x"BB";	-- JEQ @VALORATUALIZADO3 	#Se for 12, atualiza o valor e vai para a proxima configuracao
tmp(214) := CEQ & '0' & x"12";	-- CEQ @18 	#Compara com 13
tmp(215) := JEQ & '1' & x"BB";	-- JEQ @VALORATUALIZADO3 	#Se for 13, atualiza o valor e vai para a proxima configuracao
tmp(216) := CEQ & '0' & x"13";	-- CEQ @19 	#Compara com 14
tmp(217) := JEQ & '1' & x"BB";	-- JEQ @VALORATUALIZADO3 	#Se for 14, atualiza o valor e vai para a proxima configuracao
tmp(218) := CEQ & '0' & x"14";	-- CEQ @20 	#Compara com 15
tmp(219) := JEQ & '1' & x"BB";	-- JEQ @VALORATUALIZADO3 	#Se for 15, atualiza o valor e vai para a proxima configuracao
tmp(220) := NOP & '0' & x"00";	-- NOP 
tmp(221) := STA & '0' & x"0C";	-- STA @12 	#Armazena o valor das chaves no limite das unidades de milhar
tmp(222) := NOP & '0' & x"00";	-- NOP 
tmp(223) := LDI & '0' & x"80";	-- LDI $128 	# Carrega o valor 128 no acumulador
tmp(224) := STA & '1' & x"00";	-- STA @256 	# Bota o valor nos LEDS
tmp(225) := LDA & '1' & x"40";	-- LDA @320 	#Le o valor das chaves SW(7~0)
tmp(226) := CEQ & '0' & x"08";	-- CEQ @8 	#Compara com 10
tmp(227) := JEQ & '1' & x"AC";	-- JEQ @DISPLAYATUALIZADO4 	#Se for 10, atualiza o display e vai para a proxima configuracao
tmp(228) := CEQ & '0' & x"10";	-- CEQ @16 	#Compara com 11
tmp(229) := JEQ & '1' & x"AC";	-- JEQ @DISPLAYATUALIZADO4 	#Se for 11, atualiza o display e vai para a proxima configuracao
tmp(230) := CEQ & '0' & x"11";	-- CEQ @17 	#Compara com 12
tmp(231) := JEQ & '1' & x"AC";	-- JEQ @DISPLAYATUALIZADO4 	#Se for 12, atualiza o display e vai para a proxima configuracao
tmp(232) := CEQ & '0' & x"12";	-- CEQ @18 	#Compara com 13
tmp(233) := JEQ & '1' & x"AC";	-- JEQ @DISPLAYATUALIZADO4 	#Se for 13, atualiza o display e vai para a proxima configuracao
tmp(234) := CEQ & '0' & x"13";	-- CEQ @19 	#Compara com 14
tmp(235) := JEQ & '1' & x"AC";	-- JEQ @DISPLAYATUALIZADO4 	#Se for 14, atualiza o display e vai para a proxima configuracao
tmp(236) := CEQ & '0' & x"14";	-- CEQ @20 	#Compara com 15
tmp(237) := JEQ & '1' & x"AC";	-- JEQ @DISPLAYATUALIZADO4 	#Se for 15, atualiza o display e vai para a proxima configuracao
tmp(238) := NOP & '0' & x"00";	-- NOP 
tmp(239) := STA & '1' & x"24";	-- STA @292 	# Hex 4
tmp(240) := LDA & '1' & x"61";	-- LDA @353 	#Le o valor de KEY1 novamente
tmp(241) := CEQ & '0' & x"06";	-- CEQ @6 	#Compara com 0 o valor de KEY1 
tmp(242) := JEQ & '0' & x"DE";	-- JEQ @ESPERADEZENAMILHAR 	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(243) := STA & '1' & x"FE";	-- STA @510 	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(244) := LDA & '1' & x"40";	-- LDA @320 	#Le o valor das chaves SW(7~0)
tmp(245) := CEQ & '0' & x"08";	-- CEQ @8 	#Compara com 10
tmp(246) := JEQ & '1' & x"BE";	-- JEQ @VALORATUALIZADO4 	#Se for 10, atualiza o valor e vai para a proxima configuracao
tmp(247) := CEQ & '0' & x"10";	-- CEQ @16 	#Compara com 11
tmp(248) := JEQ & '1' & x"BE";	-- JEQ @VALORATUALIZADO4 	#Se for 11, atualiza o valor e vai para a proxima configuracao
tmp(249) := CEQ & '0' & x"11";	-- CEQ @17 	#Compara com 12
tmp(250) := JEQ & '1' & x"BE";	-- JEQ @VALORATUALIZADO4 	#Se for 12, atualiza o valor e vai para a proxima configuracao
tmp(251) := CEQ & '0' & x"12";	-- CEQ @18 	#Compara com 13
tmp(252) := JEQ & '1' & x"BE";	-- JEQ @VALORATUALIZADO4 	#Se for 13, atualiza o valor e vai para a proxima configuracao
tmp(253) := CEQ & '0' & x"13";	-- CEQ @19 	#Compara com 14
tmp(254) := JEQ & '1' & x"BE";	-- JEQ @VALORATUALIZADO4 	#Se for 14, atualiza o valor e vai para a proxima configuracao
tmp(255) := CEQ & '0' & x"14";	-- CEQ @20 	#Compara com 15
tmp(256) := JEQ & '1' & x"BE";	-- JEQ @VALORATUALIZADO4 	#Se for 15, atualiza o valor e vai para a proxima configuracao
tmp(257) := NOP & '0' & x"00";	-- NOP 
tmp(258) := STA & '0' & x"0D";	-- STA @13 	#Armazena o valor das chaves no limite das dezenas de milhar
tmp(259) := NOP & '0' & x"00";	-- NOP 
tmp(260) := LDA & '0' & x"06";	-- LDA @6 	#Carrega 0 no acumulador
tmp(261) := STA & '1' & x"00";	-- STA @256 	# Zera o valor nos LEDS(7~0)
tmp(262) := LDI & '0' & x"01";	-- LDI $1 	# Carrega o valor 1 no acumulador
tmp(263) := STA & '1' & x"01";	-- STA @257 	# Bota o valor nos LEDS
tmp(264) := LDA & '1' & x"40";	-- LDA @320 	#Le o valor das chaves SW(7~0)
tmp(265) := CEQ & '0' & x"08";	-- CEQ @8 	#Compara com 10
tmp(266) := JEQ & '1' & x"AF";	-- JEQ @DISPLAYATUALIZADO5 	#Se for 10, atualiza o display e vai para a proxima configuracao
tmp(267) := CEQ & '0' & x"10";	-- CEQ @16 	#Compara com 11
tmp(268) := JEQ & '1' & x"AF";	-- JEQ @DISPLAYATUALIZADO5 	#Se for 11, atualiza o display e vai para a proxima configuracao
tmp(269) := CEQ & '0' & x"11";	-- CEQ @17 	#Compara com 12
tmp(270) := JEQ & '1' & x"AF";	-- JEQ @DISPLAYATUALIZADO5 	#Se for 12, atualiza o display e vai para a proxima configuracao
tmp(271) := CEQ & '0' & x"12";	-- CEQ @18 	#Compara com 13
tmp(272) := JEQ & '1' & x"AF";	-- JEQ @DISPLAYATUALIZADO5 	#Se for 13, atualiza o display e vai para a proxima configuracao
tmp(273) := CEQ & '0' & x"13";	-- CEQ @19 	#Compara com 14
tmp(274) := JEQ & '1' & x"AF";	-- JEQ @DISPLAYATUALIZADO5 	#Se for 14, atualiza o display e vai para a proxima configuracao
tmp(275) := CEQ & '0' & x"14";	-- CEQ @20 	#Compara com 15
tmp(276) := JEQ & '1' & x"AF";	-- JEQ @DISPLAYATUALIZADO5 	#Se for 15, atualiza o display e vai para a proxima configuracao
tmp(277) := NOP & '0' & x"00";	-- NOP 
tmp(278) := STA & '1' & x"25";	-- STA @293 	# Hex 5
tmp(279) := LDA & '1' & x"61";	-- LDA @353 	#Le o valor de KEY1 novamente
tmp(280) := CEQ & '0' & x"06";	-- CEQ @6 	#Compara com 0 o valor de KEY1
tmp(281) := JEQ & '1' & x"03";	-- JEQ @ESPERACENTENAMILHAR 	#Se for igual a 0, ficar em LOOP "esperando" o valor mudar
tmp(282) := STA & '1' & x"FE";	-- STA @510 	#Se for diferente de 0, Limpa a leitura de KEY1
tmp(283) := LDA & '1' & x"40";	-- LDA @320 	#Le o valor das chaves SW(7~0)
tmp(284) := CEQ & '0' & x"08";	-- CEQ @8 	#Compara com 10
tmp(285) := JEQ & '1' & x"C1";	-- JEQ @VALORATUALIZADO5 	#Se for 10, atualiza o valor e vai para a proxima configuracao
tmp(286) := CEQ & '0' & x"10";	-- CEQ @16 	#Compara com 11
tmp(287) := JEQ & '1' & x"C1";	-- JEQ @VALORATUALIZADO5 	#Se for 11, atualiza o valor e vai para a proxima configuracao
tmp(288) := CEQ & '0' & x"11";	-- CEQ @17 	#Compara com 12
tmp(289) := JEQ & '1' & x"C1";	-- JEQ @VALORATUALIZADO5 	#Se for 12, atualiza o valor e vai para a proxima configuracao
tmp(290) := CEQ & '0' & x"12";	-- CEQ @18 	#Compara com 13
tmp(291) := JEQ & '1' & x"C1";	-- JEQ @VALORATUALIZADO5 	#Se for 13, atualiza o valor e vai para a proxima configuracao
tmp(292) := CEQ & '0' & x"13";	-- CEQ @19 	#Compara com 14
tmp(293) := JEQ & '1' & x"C1";	-- JEQ @VALORATUALIZADO5 	#Se for 14, atualiza o valor e vai para a proxima configuracao
tmp(294) := CEQ & '0' & x"14";	-- CEQ @20 	#Compara com 15
tmp(295) := JEQ & '1' & x"C1";	-- JEQ @VALORATUALIZADO5 	#Se for 15, atualiza o valor e vai para a proxima configuracao
tmp(296) := NOP & '0' & x"00";	-- NOP 
tmp(297) := STA & '0' & x"0E";	-- STA @14 	#Armazena o valor das chaves no limite das centenas de milhar
tmp(298) := RET & '0' & x"00";	-- RET 	#Retorna para o LOOP principal
tmp(299) := NOP & '0' & x"00";	-- NOP 
tmp(300) := STA & '1' & x"FF";	-- STA @511 	#Limpa a leitura de KEY1
tmp(301) := NOP & '0' & x"00";	-- NOP 
tmp(302) := LDA & '0' & x"00";	-- LDA @0 	#Carrega o valor da unidade no acumulador
tmp(303) := SOMA & '0' & x"07";	-- SOMA @7     	#Incrementa 1 na unidade
tmp(304) := CEQ & '0' & x"08";	-- CEQ @8      	#Compara unidade com 10
tmp(305) := JEQ & '1' & x"34";	-- JEQ @UNIDADEPASSOU  	#Se for igual a 10, incrementa a dezena
tmp(306) := STA & '0' & x"00";	-- STA @0 	#Se for diferente de 10, armazena o valor da unidade
tmp(307) := RET & '0' & x"00";	-- RET 	#Retorna para o LOOP principal
tmp(308) := NOP & '0' & x"00";	-- NOP 
tmp(309) := LDA & '0' & x"06";	-- LDA @6 	#Carrega 0 no acumulador
tmp(310) := STA & '0' & x"00";	-- STA @0 	#Zera a unidade
tmp(311) := LDA & '0' & x"01";	-- LDA @1 	#Carrega o valor da dezena no acumulador
tmp(312) := SOMA & '0' & x"07";	-- SOMA @7     	#Incrementa 1 na dezena 
tmp(313) := CEQ & '0' & x"08";	-- CEQ @8      	#Compara dezena com 10
tmp(314) := JEQ & '1' & x"3D";	-- JEQ @DEZENAPASSOU 	#Se for igual a 10, incrementa a centena
tmp(315) := STA & '0' & x"01";	-- STA @1 	#Se for diferente de 10, armazena o valor da dezena
tmp(316) := RET & '0' & x"00";	-- RET 	#Retorna para o LOOP principal
tmp(317) := NOP & '0' & x"00";	-- NOP 
tmp(318) := LDA & '0' & x"06";	-- LDA @6 	#Carrega 0 no acumulador
tmp(319) := STA & '0' & x"01";	-- STA @1 	#Zera a dezena
tmp(320) := LDA & '0' & x"02";	-- LDA @2 	#Carrega o valor da centena no acumulador
tmp(321) := SOMA & '0' & x"07";	-- SOMA @7     	#Incrementa 1 na centena
tmp(322) := CEQ & '0' & x"08";	-- CEQ @8      	#Compara centena com 10
tmp(323) := JEQ & '1' & x"46";	-- JEQ @CENTENAPASSOU 	#Se for igual a 10, incrementa a unidade de milhar
tmp(324) := STA & '0' & x"02";	-- STA @2 	#Se for diferente de 10, armazena o valor da centena
tmp(325) := RET & '0' & x"00";	-- RET 	#Retorna para o LOOP principal
tmp(326) := NOP & '0' & x"00";	-- NOP 
tmp(327) := LDA & '0' & x"06";	-- LDA @6 	#Carrega 0 no acumulador
tmp(328) := STA & '0' & x"02";	-- STA @2 	#Zera a centena
tmp(329) := LDA & '0' & x"03";	-- LDA @3 	#Carrega o valor da unidade de milhar no acumulador
tmp(330) := SOMA & '0' & x"07";	-- SOMA @7 	#Incrementa 1 na unidade de milhar
tmp(331) := CEQ & '0' & x"08";	-- CEQ @8  	#Compara unidade de milhar com 10
tmp(332) := JEQ & '1' & x"4F";	-- JEQ @UNIDADEMILHARPASSOU 	#Se for igual a 10, incrementa a dezena de milhar
tmp(333) := STA & '0' & x"03";	-- STA @3 	#Se for diferente de 10, armazena o valor da unidade de milhar
tmp(334) := RET & '0' & x"00";	-- RET 	#Retorna para o LOOP principal
tmp(335) := NOP & '0' & x"00";	-- NOP 
tmp(336) := LDA & '0' & x"06";	-- LDA @6 	#Carrega 0 no acumulador
tmp(337) := STA & '0' & x"03";	-- STA @3 	#Zera a unidade de milhar
tmp(338) := LDA & '0' & x"04";	-- LDA @4 	#Carrega o valor da dezena de milhar no acumulador
tmp(339) := SOMA & '0' & x"07";	-- SOMA @7 	#Incrementa 1 na dezena de milhar
tmp(340) := CEQ & '0' & x"08";	-- CEQ @8  	#Compara dezena de milhar com 10
tmp(341) := JEQ & '1' & x"58";	-- JEQ @DEZENAMILHARPASSOU 	#Se for igual a 10, incrementa a centena de milhar
tmp(342) := STA & '0' & x"04";	-- STA @4 	#Se for diferente de 10, armazena o valor da dezena de milhar
tmp(343) := RET & '0' & x"00";	-- RET 	#Retorna para o LOOP principal
tmp(344) := NOP & '0' & x"00";	-- NOP 
tmp(345) := LDA & '0' & x"06";	-- LDA @6 	#Carrega 0 no acumulador
tmp(346) := STA & '0' & x"04";	-- STA @4 	#Zera a dezena de milhar
tmp(347) := LDA & '0' & x"05";	-- LDA @5 	#Carrega o valor da centena de milhar no acumulador
tmp(348) := SOMA & '0' & x"07";	-- SOMA @7 	#Incrementa 1 na centena de milhar
tmp(349) := CEQ & '0' & x"08";	-- CEQ @8  	#Compara centena de milhar com 10
tmp(350) := JEQ & '1' & x"61";	-- JEQ @CENTENAMILHARPASSOU 	#Se for igual a 10, incrementa a unidade de milhao
tmp(351) := STA & '0' & x"05";	-- STA @5 	#Se for diferente de 10, armazena o valor da centena de milhar
tmp(352) := RET & '0' & x"00";	-- RET 	#Retorna para o LOOP principal
tmp(353) := NOP & '0' & x"00";	-- NOP 
tmp(354) := LDA & '0' & x"06";	-- LDA @6 	#Carrega 0 no acumulador
tmp(355) := STA & '0' & x"05";	-- STA @5 	#Zera a centena de milhar
tmp(356) := LDI & '0' & x"01";	-- LDI $1 	#Carrega 1 no acumulador
tmp(357) := STA & '1' & x"02";	-- STA @258 	#Acende o LED(9)
tmp(358) := STA & '0' & x"0F";	-- STA @15 	#Ativa a flag de inibir incremento
tmp(359) := RET & '0' & x"00";	-- RET 	#Retorna para o LOOP principal
tmp(360) := NOP & '0' & x"00";	-- NOP  	#Atualiza os valores dos HEX
tmp(361) := LDA & '0' & x"00";	-- LDA @0 	#Le o valor das unidades
tmp(362) := STA & '1' & x"20";	-- STA @288 	#Armazena o valor das unidades no HEX0
tmp(363) := LDA & '0' & x"01";	-- LDA @1 	#Le o valor das dezenas
tmp(364) := STA & '1' & x"21";	-- STA @289 	#Armazena o valor das dezenas no HEX1
tmp(365) := LDA & '0' & x"02";	-- LDA @2 	#Le o valor das centenas
tmp(366) := STA & '1' & x"22";	-- STA @290 	#Armazena o valor das centenas no HEX2
tmp(367) := LDA & '0' & x"03";	-- LDA @3 	#Le o valor das unidades de milhar
tmp(368) := STA & '1' & x"23";	-- STA @291 	#Armazena o valor das unidades de milhar no HEX3
tmp(369) := LDA & '0' & x"04";	-- LDA @4 	#Le o valor das dezenas de milhar
tmp(370) := STA & '1' & x"24";	-- STA @292 	#Armazena o valor das dezenas de milhar no HEX4
tmp(371) := LDA & '0' & x"05";	-- LDA @5 	#Le o valor das centenas de milhar
tmp(372) := STA & '1' & x"25";	-- STA @293 	#Armazena o valor das centenas de milhar no HEX5
tmp(373) := RET & '0' & x"00";	-- RET 	#Retorna para o LOOP principal
tmp(374) := NOP & '0' & x"00";	-- NOP 
tmp(375) := LDA & '0' & x"00";	-- LDA @0 	#Le o valor das unidades
tmp(376) := CEQ & '0' & x"09";	-- CEQ @9 	# Compara com o valor limite das unidades
tmp(377) := JEQ & '1' & x"7B";	-- JEQ @CHECADEZENA 	#Se for igual, checa se ocorre com as dezenas
tmp(378) := RET & '0' & x"00";	-- RET 	#Se for diferente, retorna para o LOOP principal
tmp(379) := NOP & '0' & x"00";	-- NOP 
tmp(380) := LDA & '0' & x"01";	-- LDA @1 	#Le o valor das dezenas
tmp(381) := CEQ & '0' & x"0A";	-- CEQ @10 	#Compara com o valor limite das dezenas
tmp(382) := JEQ & '1' & x"80";	-- JEQ @CHECACENTENA 	#Se for igual, checa se ocorre com as centenas
tmp(383) := RET & '0' & x"00";	-- RET 	#Se for diferente, retorna para o LOOP principal
tmp(384) := NOP & '0' & x"00";	-- NOP 
tmp(385) := LDA & '0' & x"02";	-- LDA @2 	#Le o valor das centenas
tmp(386) := CEQ & '0' & x"0B";	-- CEQ @11 	#Compara com o valor limite das centenas
tmp(387) := JEQ & '1' & x"85";	-- JEQ @CHECAUNIDADEMILHAR 	#Se for igual, checa se ocorre com as unidades de milhar
tmp(388) := RET & '0' & x"00";	-- RET 	#Se for diferente, retorna para o LOOP principal
tmp(389) := NOP & '0' & x"00";	-- NOP 
tmp(390) := LDA & '0' & x"03";	-- LDA @3 	# Le o valor das unidades de milhar
tmp(391) := CEQ & '0' & x"0C";	-- CEQ @12 	# Compara com o valor limite das unidades de milhar 
tmp(392) := JEQ & '1' & x"8A";	-- JEQ @CHECADEZENAMILHAR 	#Se for igual, checa se ocorre com as dezenas de milhar
tmp(393) := RET & '0' & x"00";	-- RET 	#Se for diferente, retorna para o LOOP principal
tmp(394) := NOP & '0' & x"00";	-- NOP 
tmp(395) := LDA & '0' & x"04";	-- LDA @4 	# Le o valor das dezenas de milhar
tmp(396) := CEQ & '0' & x"0D";	-- CEQ @13 	# Compara com o valor limite das dezenas de milhar 
tmp(397) := JEQ & '1' & x"8F";	-- JEQ @CHECACENTENAMILHAR 	#Se for igual, checa se ocorre com as centenas de milhar
tmp(398) := RET & '0' & x"00";	-- RET 	#Se for diferente, retorna para o LOOP principal
tmp(399) := NOP & '0' & x"00";	-- NOP 
tmp(400) := LDA & '0' & x"05";	-- LDA @5 	# Le o valor das centenas de milhar
tmp(401) := CEQ & '0' & x"0E";	-- CEQ @14 	# Compara com o valor limite das centenas de milhar 
tmp(402) := JEQ & '1' & x"94";	-- JEQ @BATEUNOLIMITE 	#Se for igual, indica que o limite foi batido
tmp(403) := RET & '0' & x"00";	-- RET 	#Se for diferente, retorna para o LOOP principal
tmp(404) := NOP & '0' & x"00";	-- NOP 
tmp(405) := LDI & '0' & x"01";	-- LDI $1 	#Atribui o valor 1 no acumulador
tmp(406) := STA & '0' & x"0F";	-- STA @15 	#Ativa a flag de parar contagem
tmp(407) := STA & '1' & x"02";	-- STA @258 	#Ativa o LED de limite atingido 
tmp(408) := RET & '0' & x"00";	-- RET 	#Retorna pro LOOP principal
tmp(409) := NOP & '0' & x"00";	-- NOP  	#Trava a contagem
tmp(410) := LDI & '0' & x"01";	-- LDI $1
tmp(411) := STA & '1' & x"00";	-- STA @256
tmp(412) := LDA & '1' & x"64";	-- LDA @356 	#Le o valor do botao FPGA
tmp(413) := CEQ & '0' & x"06";	-- CEQ @6 	#Compara com 0 o botao FPGA
tmp(414) := JEQ & '1' & x"99";	-- JEQ @TRAVA 	#Se for igual, continua travado
tmp(415) := JMP & '0' & x"00";	-- JMP @RESTART 	#Se for diferente, reinicia a contagem
tmp(416) := NOP & '0' & x"00";	-- NOP  	#Atualiza o display das unidades
tmp(417) := LDI & '0' & x"09";	-- LDI $9
tmp(418) := JMP & '0' & x"5A";	-- JMP @RETORNA 
tmp(419) := NOP & '0' & x"00";	-- NOP  	# Atualiza o display das dezenas
tmp(420) := LDI & '0' & x"09";	-- LDI $9
tmp(421) := JMP & '0' & x"7F";	-- JMP @RETORNA2
tmp(422) := NOP & '0' & x"00";	-- NOP  	# Atualiza o display das centenas
tmp(423) := LDI & '0' & x"09";	-- LDI $9
tmp(424) := JMP & '0' & x"A4";	-- JMP @RETORNA3
tmp(425) := NOP & '0' & x"00";	-- NOP  	# Atualiza o display das unidades de milhar
tmp(426) := LDI & '0' & x"09";	-- LDI $9
tmp(427) := JMP & '0' & x"C9";	-- JMP @RETORNA4
tmp(428) := NOP & '0' & x"00";	-- NOP  	# Atualiza o display das dezenas de milhar
tmp(429) := LDI & '0' & x"09";	-- LDI $9
tmp(430) := JMP & '0' & x"EE";	-- JMP @RETORNA5
tmp(431) := NOP & '0' & x"00";	-- NOP  	# Atualiza o display das centenas de milhar
tmp(432) := LDI & '0' & x"09";	-- LDI $9
tmp(433) := JMP & '1' & x"15";	-- JMP @RETORNA6
tmp(434) := NOP & '0' & x"00";	-- NOP  	# Atualiza o valor das unidades
tmp(435) := LDI & '0' & x"09";	-- LDI $9
tmp(436) := JMP & '0' & x"6D";	-- JMP @RETORNA7
tmp(437) := NOP & '0' & x"00";	-- NOP  	# Atualiza o valor das dezenas
tmp(438) := LDI & '0' & x"09";	-- LDI $9
tmp(439) := JMP & '0' & x"92";	-- JMP @RETORNA8
tmp(440) := NOP & '0' & x"00";	-- NOP  	# Atualiza o valor das centenas
tmp(441) := LDI & '0' & x"09";	-- LDI $9
tmp(442) := JMP & '0' & x"B7";	-- JMP @RETORNA9
tmp(443) := NOP & '0' & x"00";	-- NOP  	# Atualiza o valor das unidades de milhar
tmp(444) := LDI & '0' & x"09";	-- LDI $9
tmp(445) := JMP & '0' & x"DC";	-- JMP @RETORNA10
tmp(446) := NOP & '0' & x"00";	-- NOP  	# Atualiza o valor das dezenas de milhar
tmp(447) := LDI & '0' & x"09";	-- LDI $9
tmp(448) := JMP & '1' & x"01";	-- JMP @RETORNA11
tmp(449) := NOP & '0' & x"00";	-- NOP  	# Atualiza o valor das centenas de milhar
tmp(450) := LDI & '0' & x"09";	-- LDI $9
tmp(451) := JMP & '1' & x"28";	-- JMP @RETORNA12
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;